///////////////////////////////////////////////////////////////////////////////
// vim:set shiftwidth=3 softtabstop=3 expandtab:
// $Id: packer 2008-03-13 gac1 $
//
// Module: packer.v
// Project: NF2.1
// Description: defines a module for the user data path
//
///////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ps

module packer
   #(
      parameter DATA_WIDTH = 64,
      parameter CTRL_WIDTH = DATA_WIDTH/8,
      parameter UDP_REG_SRC_WIDTH = 2,
      parameter IO_QUEUE_STAGE_NUM = `IO_QUEUE_STAGE_NUM,
      parameter TIME_WIDTH = 64
   )
   (
      // --- data path interface
      output [DATA_WIDTH-1:0] 		out_data,
      output [CTRL_WIDTH-1:0] 		out_ctrl,
      output 				out_wr,
      input 				out_rdy,

      input [DATA_WIDTH-1:0] 		in_data,
      input [CTRL_WIDTH-1:0] 		in_ctrl,
      input 				in_wr,
      output 				in_rdy,


      // --- Register interface
      input 				reg_req_in,
      input 				reg_ack_in,
      input 				reg_rd_wr_L_in,
      input [`UDP_REG_ADDR_WIDTH-1:0] 	reg_addr_in,
      input [`CPCI_NF2_DATA_WIDTH-1:0] 	reg_data_in,
      input [UDP_REG_SRC_WIDTH-1:0] 	reg_src_in,

      output 				reg_req_out,
      output 				reg_ack_out,
      output 				reg_rd_wr_L_out,
      output [`UDP_REG_ADDR_WIDTH-1:0] 	reg_addr_out,
      output [`CPCI_NF2_DATA_WIDTH-1:0] reg_data_out,
      output [UDP_REG_SRC_WIDTH-1:0] 	reg_src_out,

      // misc
      input 				clk,
      input 				reset
   );

   // Include the log2 function
   `LOG2_FUNC

   //------------------------- Signals-------------------------------

   wire [DATA_WIDTH-1:0]         in_fifo_data;
   wire [CTRL_WIDTH-1:0]         in_fifo_ctrl;

   reg  [DATA_WIDTH-1:0] 	 __out_data;
   reg  [CTRL_WIDTH-1:0]         old_ctrl;

   wire                          in_fifo_nearly_full;
   wire                          in_fifo_empty;

   reg                           in_fifo_rd_en;
   reg                           out_wr_int;

   wire [31:0] 			 value;

   //------------------------- Local assignments -------------------------------

   assign in_rdy     = !in_fifo_nearly_full;
   assign out_wr     = out_wr_int;
   assign out_ctrl   = in_fifo_ctrl;
   assign out_data   = __out_data;


   //------------------------- Modules-------------------------------

   fallthrough_small_fifo #(
      .WIDTH(CTRL_WIDTH+DATA_WIDTH),
      .MAX_DEPTH_BITS(2)
   ) input_fifo (
      .din           ({in_ctrl, in_data}),   // Data in
      .wr_en         (in_wr),                // Write enable
      .rd_en         (in_fifo_rd_en),        // Read the next word
      .dout          ({in_fifo_ctrl, in_fifo_data}),
      .full          (),
      .nearly_full   (in_fifo_nearly_full),
      .prog_full     (),
      .empty         (in_fifo_empty),
      .reset         (reset),
      .clk           (clk)
   );

   generic_regs
   #(
      .UDP_REG_SRC_WIDTH   (UDP_REG_SRC_WIDTH),
      .TAG                 (`PACKER_BLOCK_ADDR), // Tag -- eg. MODULE_TAG
      .REG_ADDR_WIDTH      (`PACKER_REG_ADDR_WIDTH),                 // Width of block addresses -- eg. MODULE_REG_ADDR_WIDTH
      .NUM_COUNTERS        (0),                 // Number of counters
      .NUM_SOFTWARE_REGS   (1),                 // Number of sw regs
      .NUM_HARDWARE_REGS   (0)                  // Number of hw regs
   ) packer_regs (
      .reg_req_in       (reg_req_in),
      .reg_ack_in       (reg_ack_in),
      .reg_rd_wr_L_in   (reg_rd_wr_L_in),
      .reg_addr_in      (reg_addr_in),
      .reg_data_in      (reg_data_in),
      .reg_src_in       (reg_src_in),

      .reg_req_out      (reg_req_out),
      .reg_ack_out      (reg_ack_out),
      .reg_rd_wr_L_out  (reg_rd_wr_L_out),
      .reg_addr_out     (reg_addr_out),
      .reg_data_out     (reg_data_out),
      .reg_src_out      (reg_src_out),

      // --- counters interface
      .counter_updates  (),
      .counter_decrement(),

      // --- SW regs interface
      .software_regs    (value),

      // --- HW regs interface
      .hardware_regs    (),

      .clk              (clk),
      .reset            (reset)
    );

   //------------------------- Logic-------------------------------
   /* pkt is from the cpu if it comes in on an odd numbered port */
   assign pkt_is_from_cpu = in_data[`IOQ_SRC_PORT_POS];

   always @(*) begin
      // Default values
      out_wr_int    = 0;
      in_fifo_rd_en = 0;

      if (!in_fifo_empty && out_rdy) begin
         out_wr_int    = 1;
         in_fifo_rd_en = 1;
      end

      __out_data = in_fifo_data;
      if (in_fifo_ctrl == 0) begin
	 __out_data[63:32] = value;
      end
   end

   always @(posedge clk) begin
      old_ctrl <= in_fifo_ctrl;
   end

endmodule
